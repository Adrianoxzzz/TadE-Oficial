library ieee ;
    use ieee.std_logic_1164.all ;
    use ieee.std_logic_arith.all ;
    use ieee.std_logic_unsigned.all;

entity M25P16 is
  port (
    clk
    rst
    cs
    wr
    r
  ) ;
end M25P16 ; 

architecture arch of M25P16 is

begin

end architecture ;